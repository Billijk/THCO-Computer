module vga_rom(
	input wire[6:0] ch,
	input wire[9:0] pos,
	output reg mask
);


always @(*) begin
	case(ch[6:0])
		100: begin
			case(pos[9:0])
				89, 90, 91, 92, 93, 94, 95, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 194, 195, 196, 204, 205, 206, 207, 229, 230, 231, 242, 243, 265, 266, 278, 279, 301, 302, 314, 315, 337, 338, 349, 350, 373, 374, 384, 385, 386, 409, 410, 419, 420, 421, 439, 440, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 475, 476, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 511, 512, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		101: begin
			case(pos[9:0])
				89, 90, 91, 92, 93, 94, 95, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 194, 195, 196, 199, 200, 204, 205, 206, 229, 230, 231, 235, 236, 241, 242, 243, 265, 266, 271, 272, 278, 279, 301, 302, 307, 308, 314, 315, 337, 338, 343, 344, 350, 351, 373, 374, 375, 379, 380, 386, 387, 410, 411, 412, 415, 416, 422, 423, 446, 447, 448, 449, 450, 451, 452, 458, 459, 483, 484, 485, 486, 487, 488, 493, 494, 521, 522, 523, 524:
					mask = 1;
				default: mask = 0;
			endcase
		end
		102: begin
			case(pos[9:0])
				51, 52, 87, 88, 123, 124, 159, 160, 195, 196, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 331, 332, 333, 339, 340, 367, 368, 375, 376, 403, 404, 411, 412, 439, 440, 447, 448, 475, 476, 483, 484, 511, 512, 519, 520, 547, 548:
					mask = 1;
				default: mask = 0;
			endcase
		end
		103: begin
			case(pos[9:0])
				65, 66, 67, 88, 89, 90, 91, 94, 95, 96, 97, 99, 100, 101, 102, 103, 104, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 175, 176, 177, 193, 194, 195, 200, 201, 202, 205, 206, 207, 212, 213, 229, 230, 237, 238, 242, 243, 248, 249, 265, 266, 273, 274, 278, 279, 284, 285, 301, 302, 309, 310, 314, 315, 320, 321, 337, 338, 345, 346, 350, 351, 356, 357, 373, 374, 375, 380, 381, 382, 386, 387, 392, 393, 409, 410, 411, 412, 413, 414, 415, 416, 417, 422, 423, 424, 427, 428, 445, 446, 447, 448, 449, 450, 451, 452, 458, 459, 460, 461, 462, 463, 464, 481, 482, 484, 485, 486, 487, 495, 496, 497, 498, 499, 517, 518, 532, 533, 534, 553, 554:
					mask = 1;
				default: mask = 0;
			endcase
		end
		104: begin
			case(pos[9:0])
				79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 195, 196, 230, 231, 265, 266, 301, 302, 337, 338, 373, 374, 375, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495:
					mask = 1;
				default: mask = 0;
			endcase
		end
		105: begin
			case(pos[9:0])
				121, 122, 134, 135, 157, 158, 170, 171, 193, 194, 206, 207, 229, 230, 242, 243, 260, 261, 265, 266, 278, 279, 295, 296, 297, 298, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 331, 332, 333, 334, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 368, 369, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 422, 423, 458, 459, 494, 495, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		106: begin
			case(pos[9:0])
				103, 104, 121, 122, 140, 141, 157, 158, 176, 177, 193, 194, 212, 213, 229, 230, 248, 249, 265, 266, 284, 285, 301, 302, 319, 320, 321, 332, 333, 337, 338, 354, 355, 356, 367, 368, 369, 370, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 403, 404, 405, 406, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 440, 441, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461:
					mask = 1;
				default: mask = 0;
			endcase
		end
		107: begin
			case(pos[9:0])
				115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 235, 236, 270, 271, 272, 273, 305, 306, 307, 308, 309, 310, 340, 341, 342, 345, 346, 347, 348, 375, 376, 377, 382, 383, 384, 385, 410, 411, 412, 419, 420, 421, 422, 445, 446, 447, 456, 457, 458, 459, 481, 482, 493, 494, 495, 517, 530, 531, 567:
					mask = 1;
				default: mask = 0;
			endcase
		end
		108: begin
			case(pos[9:0])
				115, 116, 134, 135, 151, 152, 170, 171, 187, 188, 206, 207, 223, 224, 242, 243, 259, 260, 278, 279, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 422, 423, 458, 459, 494, 495, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		109: begin
			case(pos[9:0])
				49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 158, 159, 160, 193, 194, 229, 230, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 374, 375, 376, 409, 410, 445, 446, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563, 564, 565, 566, 567:
					mask = 1;
				default: mask = 0;
			endcase
		end
		110: begin
			case(pos[9:0])
				85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 195, 196, 230, 231, 265, 266, 301, 302, 337, 338, 373, 374, 375, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495:
					mask = 1;
				default: mask = 0;
			endcase
		end
		111: begin
			case(pos[9:0])
				53, 54, 55, 56, 57, 58, 59, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 158, 159, 160, 161, 168, 169, 170, 193, 194, 195, 205, 206, 207, 229, 230, 242, 243, 265, 266, 278, 279, 301, 302, 314, 315, 337, 338, 350, 351, 373, 374, 375, 385, 386, 387, 410, 411, 412, 419, 420, 421, 422, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 521, 522, 523, 524, 525, 526, 527:
					mask = 1;
				default: mask = 0;
			endcase
		end
		112: begin
			case(pos[9:0])
				85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 100, 101, 102, 103, 104, 105, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 136, 137, 138, 139, 140, 141, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 195, 196, 206, 207, 230, 231, 242, 243, 265, 266, 267, 278, 279, 301, 302, 314, 315, 337, 338, 350, 351, 373, 374, 385, 386, 387, 409, 410, 411, 412, 419, 420, 421, 422, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 521, 522, 523, 524, 525, 526, 527:
					mask = 1;
				default: mask = 0;
			endcase
		end
		113: begin
			case(pos[9:0])
				90, 91, 92, 93, 94, 95, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 194, 195, 196, 204, 205, 206, 207, 229, 230, 231, 242, 243, 265, 266, 278, 279, 301, 302, 314, 315, 337, 338, 349, 350, 373, 374, 384, 385, 386, 409, 410, 419, 420, 421, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 460, 461, 462, 463, 464, 465, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 496, 497, 498, 499, 500, 501, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 532, 533, 534, 535, 536, 537:
					mask = 1;
				default: mask = 0;
			endcase
		end
		114: begin
			case(pos[9:0])
				121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 231, 232, 233, 266, 267, 268, 302, 303, 337, 338, 373, 374, 409, 410, 445, 446, 447, 481, 482, 483, 484, 485, 486, 518, 519, 520, 521, 522, 556, 557, 558:
					mask = 1;
				default: mask = 0;
			endcase
		end
		115: begin
			case(pos[9:0])
				123, 124, 125, 126, 133, 134, 158, 159, 160, 161, 162, 163, 169, 170, 171, 194, 195, 196, 197, 198, 199, 200, 206, 207, 229, 230, 231, 234, 235, 236, 242, 243, 265, 266, 271, 272, 278, 279, 301, 302, 307, 308, 309, 314, 315, 337, 338, 343, 344, 345, 350, 351, 373, 374, 380, 381, 386, 387, 409, 410, 416, 417, 418, 421, 422, 423, 445, 446, 452, 453, 454, 455, 456, 457, 458, 482, 483, 489, 490, 491, 492, 493, 494, 526, 527, 528, 529:
					mask = 1;
				default: mask = 0;
			endcase
		end
		116: begin
			case(pos[9:0])
				49, 50, 85, 86, 121, 122, 157, 158, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 301, 302, 313, 314, 315, 337, 338, 350, 351, 373, 374, 386, 387, 409, 410, 422, 423, 445, 446, 458, 459, 481, 482, 494, 495:
					mask = 1;
				default: mask = 0;
			endcase
		end
		117: begin
			case(pos[9:0])
				85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 205, 206, 207, 242, 243, 278, 279, 314, 315, 349, 350, 384, 385, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495:
					mask = 1;
				default: mask = 0;
			endcase
		end
		118: begin
			case(pos[9:0])
				85, 86, 87, 121, 122, 123, 124, 125, 157, 158, 159, 160, 161, 162, 163, 164, 196, 197, 198, 199, 200, 201, 202, 203, 236, 237, 238, 239, 240, 241, 242, 275, 276, 277, 278, 279, 314, 315, 347, 348, 349, 350, 351, 380, 381, 382, 383, 384, 385, 413, 414, 415, 416, 417, 418, 419, 446, 447, 448, 449, 450, 451, 452, 481, 482, 483, 484, 485, 517, 518, 519:
					mask = 1;
				default: mask = 0;
			endcase
		end
		119: begin
			case(pos[9:0])
				49, 50, 51, 52, 53, 54, 55, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 170, 171, 203, 204, 205, 206, 207, 236, 237, 238, 239, 240, 241, 269, 270, 271, 272, 273, 274, 305, 306, 307, 341, 342, 343, 344, 345, 346, 380, 381, 382, 383, 384, 385, 419, 420, 421, 422, 423, 457, 458, 459, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 553, 554, 555, 556, 557, 558, 559:
					mask = 1;
				default: mask = 0;
			endcase
		end
		120: begin
			case(pos[9:0])
				49, 63, 85, 86, 98, 99, 121, 122, 123, 133, 134, 135, 157, 158, 159, 160, 161, 167, 168, 169, 170, 171, 195, 196, 197, 198, 202, 203, 204, 205, 232, 233, 234, 235, 236, 237, 238, 239, 240, 269, 270, 271, 272, 273, 274, 306, 307, 308, 309, 340, 341, 342, 343, 344, 345, 346, 347, 375, 376, 377, 378, 381, 382, 383, 384, 410, 411, 412, 413, 418, 419, 420, 421, 445, 446, 447, 456, 457, 458, 459, 481, 482, 493, 494, 495, 517, 530, 531, 567:
					mask = 1;
				default: mask = 0;
			endcase
		end
		121: begin
			case(pos[9:0])
				68, 69, 85, 86, 87, 104, 105, 121, 122, 123, 124, 125, 140, 141, 157, 158, 159, 160, 161, 162, 163, 164, 176, 177, 196, 197, 198, 199, 200, 201, 202, 203, 211, 212, 235, 236, 237, 238, 239, 240, 241, 242, 245, 246, 247, 248, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 313, 314, 315, 316, 317, 346, 347, 348, 349, 350, 351, 379, 380, 381, 382, 383, 384, 385, 413, 414, 415, 416, 417, 418, 446, 447, 448, 449, 450, 451, 452, 481, 482, 483, 484, 485, 517, 518, 519:
					mask = 1;
				default: mask = 0;
			endcase
		end
		122: begin
			case(pos[9:0])
				85, 86, 98, 99, 121, 122, 133, 134, 135, 157, 158, 167, 168, 169, 170, 171, 193, 194, 202, 203, 204, 205, 206, 207, 229, 230, 236, 237, 238, 239, 242, 243, 265, 266, 271, 272, 273, 274, 278, 279, 301, 302, 305, 306, 307, 308, 314, 315, 337, 338, 340, 341, 342, 343, 350, 351, 373, 374, 375, 376, 377, 386, 387, 409, 410, 411, 412, 422, 423, 445, 446, 458, 459:
					mask = 1;
				default: mask = 0;
			endcase
		end
		123: begin
			case(pos[9:0])
				91, 92, 127, 128, 163, 164, 198, 199, 200, 201, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 331, 332, 333, 355, 356, 357, 367, 368, 392, 393, 403, 404, 428, 429, 439, 440, 464, 465:
					mask = 1;
				default: mask = 0;
			endcase
		end
		124: begin
			case(pos[9:0])
				256, 257, 258, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 285, 292, 293, 294, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 321, 328, 329, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357:
					mask = 1;
				default: mask = 0;
			endcase
		end
		125: begin
			case(pos[9:0])
				115, 116, 140, 141, 151, 152, 176, 177, 187, 188, 212, 213, 223, 224, 225, 247, 248, 249, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 274, 275, 276, 277, 278, 279, 280, 281, 282, 283, 284, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 309, 310, 311, 312, 313, 314, 315, 316, 317, 318, 319, 320, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 378, 379, 380, 381, 415, 416, 451, 452, 487, 488:
					mask = 1;
				default: mask = 0;
			endcase
		end
		126: begin
			case(pos[9:0])
				55, 56, 57, 90, 91, 92, 93, 125, 126, 127, 128, 129, 161, 162, 163, 197, 198, 233, 234, 270, 271, 307, 308, 344, 345, 381, 382, 417, 418, 452, 453, 454, 486, 487, 488, 489, 490, 522, 523, 524, 525, 558, 559, 560:
					mask = 1;
				default: mask = 0;
			endcase
		end
		32: begin
			mask = 0;
		end
		33: begin
			case(pos[9:0])
				223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 241, 242, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 276, 277, 278, 279, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 312, 313, 314, 315, 349, 350:
					mask = 1;
				default: mask = 0;
			endcase
		end
		34: begin
			case(pos[9:0])
				115, 116, 117, 118, 119, 120, 121, 151, 152, 153, 154, 155, 156, 157, 187, 188, 189, 190, 191, 192, 193, 223, 224, 225, 226, 227, 228, 229, 331, 332, 333, 334, 335, 336, 337, 367, 368, 369, 370, 371, 372, 373, 403, 404, 405, 406, 407, 408, 409, 439, 440, 441, 442, 443, 444, 445:
					mask = 1;
				default: mask = 0;
			endcase
		end
		35: begin
			case(pos[9:0])
				57, 58, 86, 87, 93, 94, 122, 123, 129, 130, 158, 159, 165, 166, 168, 169, 170, 171, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 273, 274, 302, 303, 309, 310, 312, 313, 314, 315, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 441, 442, 443, 444, 445, 446, 447, 453, 454, 482, 483, 489, 490, 518, 519, 525, 526, 554, 555:
					mask = 1;
				default: mask = 0;
			endcase
		end
		36: begin
			case(pos[9:0])
				84, 85, 86, 87, 97, 98, 119, 120, 121, 122, 123, 124, 134, 154, 155, 156, 157, 158, 159, 160, 161, 170, 171, 190, 191, 195, 196, 197, 206, 207, 225, 226, 232, 233, 234, 241, 242, 243, 244, 245, 246, 261, 262, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 280, 281, 282, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 330, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 350, 351, 366, 367, 368, 369, 370, 371, 378, 379, 380, 386, 387, 405, 406, 414, 415, 416, 421, 422, 441, 442, 451, 452, 453, 454, 455, 456, 457, 458, 478, 479, 487, 488, 489, 490, 491, 492, 493, 525, 526, 527, 528:
					mask = 1;
				default: mask = 0;
			endcase
		end
		37: begin
			case(pos[9:0])
				27, 45, 46, 47, 48, 49, 62, 63, 80, 81, 82, 83, 84, 85, 86, 96, 97, 98, 99, 115, 116, 117, 118, 119, 120, 121, 122, 123, 131, 132, 133, 151, 152, 153, 158, 159, 165, 166, 167, 168, 187, 188, 194, 195, 200, 201, 202, 223, 224, 229, 230, 231, 234, 235, 236, 237, 259, 260, 261, 262, 263, 264, 265, 266, 267, 269, 270, 271, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 309, 310, 311, 312, 313, 333, 334, 335, 336, 337, 338, 339, 340, 344, 345, 346, 347, 348, 349, 350, 372, 373, 374, 375, 379, 380, 381, 382, 383, 384, 385, 386, 387, 407, 408, 409, 415, 416, 417, 422, 423, 441, 442, 443, 444, 451, 452, 458, 459, 476, 477, 478, 487, 488, 493, 494, 495, 511, 512, 513, 523, 524, 525, 526, 527, 528, 529, 530, 531, 547, 560, 561, 562, 563, 564, 565, 566:
					mask = 1;
				default: mask = 0;
			endcase
		end
		38: begin
			case(pos[9:0])
				56, 57, 58, 59, 60, 91, 92, 93, 94, 95, 96, 97, 118, 119, 120, 121, 122, 126, 127, 128, 129, 130, 131, 132, 133, 134, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 168, 169, 170, 171, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 205, 206, 207, 223, 224, 225, 230, 231, 232, 233, 234, 242, 243, 259, 260, 267, 268, 269, 270, 271, 278, 279, 295, 296, 303, 304, 305, 306, 307, 308, 314, 315, 331, 332, 333, 338, 339, 340, 342, 343, 344, 345, 350, 351, 367, 368, 369, 370, 371, 372, 373, 374, 375, 380, 381, 382, 385, 386, 387, 404, 405, 406, 407, 408, 409, 410, 417, 418, 419, 421, 422, 441, 442, 443, 444, 445, 454, 455, 456, 457, 458, 486, 487, 488, 489, 490, 491, 492, 493, 494, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 558, 559, 560, 561, 565, 566, 567:
					mask = 1;
				default: mask = 0;
			endcase
		end
		39: begin
			case(pos[9:0])
				259, 260, 261, 262, 263, 264, 265, 295, 296, 297, 298, 299, 300, 301, 331, 332, 333, 334, 335, 336, 337, 367, 368, 369, 370, 371, 372, 373:
					mask = 1;
				default: mask = 0;
			endcase
		end
		40: begin
			case(pos[9:0])
				160, 161, 162, 163, 164, 165, 166, 167, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 262, 263, 264, 265, 266, 267, 276, 277, 278, 279, 280, 281, 297, 298, 299, 300, 314, 315, 316, 317, 318, 332, 333, 334, 335, 352, 353, 354, 355, 367, 368, 369, 390, 391, 392, 402, 403, 404, 427, 428, 429, 439, 464:
					mask = 1;
				default: mask = 0;
			endcase
		end
		41: begin
			case(pos[9:0])
				115, 140, 150, 151, 152, 175, 176, 177, 187, 188, 189, 210, 211, 212, 224, 225, 226, 227, 244, 245, 246, 247, 261, 262, 263, 264, 279, 280, 281, 282, 298, 299, 300, 301, 302, 303, 312, 313, 314, 315, 316, 317, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 412, 413, 414, 415, 416, 417, 418, 419:
					mask = 1;
				default: mask = 0;
			endcase
		end
		42: begin
			case(pos[9:0])
				82, 87, 117, 118, 123, 124, 154, 155, 158, 159, 191, 194, 227, 228, 229, 230, 259, 260, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 295, 296, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 335, 336, 337, 338, 371, 374, 406, 407, 410, 411, 441, 442, 443, 447, 448, 478, 483:
					mask = 1;
				default: mask = 0;
			endcase
		end
		43: begin
			case(pos[9:0])
				55, 56, 91, 92, 127, 128, 163, 164, 199, 200, 235, 236, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 379, 380, 415, 416, 451, 452, 487, 488, 523, 524, 559, 560:
					mask = 1;
				default: mask = 0;
			endcase
		end
		44: begin
			case(pos[9:0])
				175, 176, 211, 212, 240, 241, 242, 246, 247, 248, 275, 276, 277, 278, 279, 280, 281, 282, 283, 311, 312, 313, 314, 315, 316, 317, 318, 319, 347, 348, 349, 350, 351, 352, 353, 354, 384, 385, 386, 387, 388:
					mask = 1;
				default: mask = 0;
			endcase
		end
		45: begin
			case(pos[9:0])
				163, 164, 199, 200, 235, 236, 271, 272, 307, 308, 343, 344, 379, 380, 415, 416, 451, 452:
					mask = 1;
				default: mask = 0;
			endcase
		end
		46: begin
			case(pos[9:0])
				240, 241, 242, 275, 276, 277, 278, 279, 311, 312, 313, 314, 315, 347, 348, 349, 350, 351, 384, 385, 386:
					mask = 1;
				default: mask = 0;
			endcase
		end
		47: begin
			case(pos[9:0])
				102, 135, 136, 137, 138, 169, 170, 171, 172, 173, 174, 203, 204, 205, 206, 207, 236, 237, 238, 239, 240, 241, 270, 271, 272, 273, 274, 275, 303, 304, 305, 306, 307, 308, 337, 338, 339, 340, 341, 342, 371, 372, 373, 374, 375, 404, 405, 406, 407, 408, 409, 439, 440, 441, 442, 443, 475, 476:
					mask = 1;
				default: mask = 0;
			endcase
		end
		48: begin
			case(pos[9:0])
				50, 51, 52, 53, 54, 55, 56, 57, 58, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 154, 155, 156, 157, 165, 166, 167, 168, 169, 170, 189, 190, 191, 200, 201, 205, 206, 207, 225, 226, 235, 236, 242, 243, 261, 262, 270, 271, 278, 279, 297, 298, 305, 306, 314, 315, 333, 334, 340, 341, 350, 351, 369, 370, 371, 375, 376, 385, 386, 387, 406, 407, 408, 409, 410, 411, 419, 420, 421, 422, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 518, 519, 520, 521, 522, 523, 524, 525, 526:
					mask = 1;
				default: mask = 0;
			endcase
		end
		49: begin
			case(pos[9:0])
				84, 119, 120, 121, 134, 135, 155, 156, 170, 171, 190, 191, 192, 206, 207, 226, 227, 242, 243, 261, 262, 278, 279, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 422, 423, 458, 459, 494, 495, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		50: begin
			case(pos[9:0])
				83, 98, 99, 118, 119, 120, 133, 134, 135, 154, 155, 168, 169, 170, 171, 189, 190, 203, 204, 205, 206, 207, 225, 226, 238, 239, 240, 242, 243, 261, 262, 273, 274, 275, 278, 279, 297, 298, 308, 309, 310, 314, 315, 333, 334, 342, 343, 344, 345, 350, 351, 369, 370, 371, 372, 377, 378, 379, 380, 386, 387, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 422, 423, 443, 444, 445, 446, 447, 448, 449, 450, 458, 459, 480, 481, 482, 483, 484, 494, 495, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		51: begin
			case(pos[9:0])
				98, 99, 118, 119, 134, 135, 153, 154, 161, 162, 170, 171, 189, 190, 197, 198, 206, 207, 225, 226, 233, 234, 242, 243, 261, 262, 269, 270, 278, 279, 297, 298, 304, 305, 306, 314, 315, 333, 334, 335, 340, 341, 342, 343, 349, 350, 370, 371, 372, 373, 374, 375, 376, 378, 379, 380, 384, 385, 386, 406, 407, 408, 409, 410, 411, 412, 414, 415, 416, 417, 418, 419, 420, 421, 422, 443, 444, 445, 446, 447, 451, 452, 453, 454, 455, 456, 457, 488, 489, 490, 491:
					mask = 1;
				default: mask = 0;
			endcase
		end
		52: begin
			case(pos[9:0])
				57, 58, 59, 92, 93, 94, 95, 126, 127, 128, 129, 130, 131, 160, 161, 162, 163, 166, 167, 195, 196, 197, 198, 202, 203, 229, 230, 231, 232, 238, 239, 263, 264, 265, 266, 267, 274, 275, 298, 299, 300, 301, 310, 311, 333, 334, 335, 346, 347, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 490, 491, 526, 527, 562, 563:
					mask = 1;
				default: mask = 0;
			endcase
		end
		53: begin
			case(pos[9:0])
				117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 170, 171, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 206, 207, 225, 226, 233, 234, 242, 243, 261, 262, 269, 270, 278, 279, 297, 298, 305, 306, 314, 315, 333, 334, 341, 342, 350, 351, 369, 370, 377, 378, 379, 385, 386, 405, 406, 414, 415, 416, 420, 421, 422, 441, 442, 450, 451, 452, 453, 454, 455, 456, 457, 477, 478, 487, 488, 489, 490, 491, 492, 493, 524, 525, 526, 527:
					mask = 1;
				default: mask = 0;
			endcase
		end
		54: begin
			case(pos[9:0])
				87, 88, 89, 90, 91, 92, 93, 94, 95, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 191, 192, 193, 194, 197, 198, 203, 204, 205, 206, 226, 227, 228, 232, 233, 241, 242, 243, 262, 263, 268, 269, 278, 279, 297, 298, 299, 304, 305, 314, 315, 333, 334, 340, 341, 350, 351, 369, 370, 376, 377, 386, 387, 405, 406, 412, 413, 414, 421, 422, 423, 441, 442, 448, 449, 450, 451, 456, 457, 458, 477, 478, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 522, 523, 524, 525, 526, 527, 528, 529, 559, 560, 561, 562, 563:
					mask = 1;
				default: mask = 0;
			endcase
		end
		55: begin
			case(pos[9:0])
				81, 82, 117, 118, 153, 154, 171, 189, 190, 205, 206, 207, 225, 226, 239, 240, 241, 242, 243, 261, 262, 273, 274, 275, 276, 277, 278, 297, 298, 307, 308, 309, 310, 311, 312, 333, 334, 341, 342, 343, 344, 345, 346, 369, 370, 375, 376, 377, 378, 379, 405, 406, 409, 410, 411, 412, 413, 441, 442, 443, 444, 445, 446, 447, 477, 478, 479, 480, 481, 513, 514, 515:
					mask = 1;
				default: mask = 0;
			endcase
		end
		56: begin
			case(pos[9:0])
				84, 85, 86, 93, 94, 95, 96, 119, 120, 121, 122, 123, 124, 128, 129, 130, 131, 132, 133, 134, 154, 155, 156, 157, 158, 159, 160, 163, 164, 165, 166, 167, 168, 169, 170, 189, 190, 191, 195, 196, 197, 198, 199, 200, 205, 206, 207, 225, 226, 232, 233, 234, 235, 242, 243, 261, 262, 268, 269, 270, 278, 279, 297, 298, 305, 306, 314, 315, 333, 334, 341, 342, 343, 350, 351, 369, 370, 376, 377, 378, 379, 386, 387, 405, 406, 407, 411, 412, 413, 414, 415, 416, 417, 421, 422, 423, 442, 443, 444, 445, 446, 447, 448, 451, 452, 453, 454, 455, 456, 457, 458, 478, 479, 480, 481, 482, 483, 488, 489, 490, 491, 492, 493, 515, 516, 517, 518, 525, 526, 527, 528:
					mask = 1;
				default: mask = 0;
			endcase
		end
		57: begin
			case(pos[9:0])
				49, 50, 51, 52, 53, 83, 84, 85, 86, 87, 88, 89, 90, 98, 99, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 134, 135, 154, 155, 156, 161, 162, 163, 164, 170, 171, 189, 190, 191, 198, 199, 200, 206, 207, 225, 226, 235, 236, 242, 243, 261, 262, 271, 272, 278, 279, 297, 298, 307, 308, 313, 314, 333, 334, 343, 344, 349, 350, 369, 370, 371, 379, 380, 384, 385, 386, 406, 407, 408, 409, 414, 415, 418, 419, 420, 421, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 518, 519, 520, 521, 522, 523, 524, 525:
					mask = 1;
				default: mask = 0;
			endcase
		end
		58: begin
			case(pos[9:0])
				230, 231, 232, 240, 241, 242, 265, 266, 267, 268, 269, 275, 276, 277, 278, 279, 301, 302, 303, 304, 305, 311, 312, 313, 314, 315, 338, 339, 340, 348, 349, 350:
					mask = 1;
				default: mask = 0;
			endcase
		end
		59: begin
			case(pos[9:0])
				175, 176, 211, 212, 230, 231, 232, 240, 241, 242, 246, 247, 248, 265, 266, 267, 268, 269, 275, 276, 277, 278, 279, 280, 281, 282, 283, 301, 302, 303, 304, 305, 311, 312, 313, 314, 315, 316, 317, 318, 319, 338, 339, 340, 347, 348, 349, 350, 351, 352, 353, 354, 384, 385, 386, 387, 388:
					mask = 1;
				default: mask = 0;
			endcase
		end
		60: begin
			case(pos[9:0])
				127, 128, 162, 163, 164, 165, 197, 198, 199, 200, 201, 202, 232, 233, 234, 235, 236, 237, 238, 239, 267, 268, 269, 270, 273, 274, 275, 276, 303, 304, 305, 310, 311, 312, 338, 339, 340, 347, 348, 349, 373, 374, 375, 384, 385, 386, 408, 409, 410, 421, 422, 423, 445, 458:
					mask = 1;
				default: mask = 0;
			endcase
		end
		61: begin
			case(pos[9:0])
				89, 90, 94, 95, 125, 126, 130, 131, 161, 162, 166, 167, 197, 198, 202, 203, 233, 234, 238, 239, 269, 270, 274, 275, 305, 306, 310, 311, 341, 342, 346, 347, 377, 378, 382, 383, 413, 414, 418, 419, 449, 450, 454, 455, 485, 486, 490, 491, 521, 522, 526, 527:
					mask = 1;
				default: mask = 0;
			endcase
		end
		62: begin
			case(pos[9:0])
				121, 134, 156, 157, 158, 169, 170, 171, 193, 194, 195, 204, 205, 206, 230, 231, 232, 239, 240, 241, 267, 268, 269, 274, 275, 276, 303, 304, 305, 306, 309, 310, 311, 312, 340, 341, 342, 343, 344, 345, 346, 347, 377, 378, 379, 380, 381, 382, 414, 415, 416, 417, 451, 452:
					mask = 1;
				default: mask = 0;
			endcase
		end
		63: begin
			case(pos[9:0])
				151, 152, 187, 188, 205, 206, 223, 224, 232, 233, 234, 235, 236, 237, 240, 241, 242, 243, 259, 260, 261, 268, 269, 270, 271, 272, 273, 276, 277, 278, 279, 296, 297, 304, 305, 306, 307, 308, 309, 313, 314, 332, 333, 334, 339, 340, 341, 369, 370, 371, 372, 373, 374, 375, 376, 377, 406, 407, 408, 409, 410, 411, 412, 443, 444, 445, 446, 447:
					mask = 1;
				default: mask = 0;
			endcase
		end
		64: begin
			case(pos[9:0])
				17, 18, 19, 20, 21, 22, 23, 24, 25, 26, 27, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 64, 65, 66, 84, 85, 86, 87, 88, 89, 99, 100, 101, 102, 103, 118, 119, 120, 121, 138, 139, 140, 153, 154, 155, 163, 164, 165, 166, 167, 168, 169, 175, 176, 177, 188, 189, 190, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 212, 213, 224, 225, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 248, 249, 259, 260, 266, 267, 268, 269, 277, 278, 284, 285, 295, 296, 302, 303, 312, 313, 320, 321, 331, 332, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 356, 357, 367, 368, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 392, 393, 403, 404, 405, 410, 411, 412, 413, 421, 422, 427, 428, 440, 441, 442, 457, 458, 477, 478, 479, 480, 491, 492, 493, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562:
					mask = 1;
				default: mask = 0;
			endcase
		end
		65: begin
			case(pos[9:0])
				61, 62, 63, 94, 95, 96, 97, 98, 99, 127, 128, 129, 130, 131, 132, 133, 134, 160, 161, 162, 163, 164, 165, 166, 167, 193, 194, 195, 196, 197, 198, 199, 200, 202, 203, 226, 227, 228, 229, 230, 231, 232, 238, 239, 261, 262, 263, 264, 265, 274, 275, 297, 298, 310, 311, 333, 334, 335, 336, 337, 346, 347, 369, 370, 371, 372, 373, 374, 375, 376, 382, 383, 408, 409, 410, 411, 412, 413, 414, 415, 416, 418, 419, 448, 449, 450, 451, 452, 453, 454, 455, 487, 488, 489, 490, 491, 492, 493, 494, 526, 527, 528, 529, 530, 531, 565, 566, 567:
					mask = 1;
				default: mask = 0;
			endcase
		end
		66: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 197, 198, 206, 207, 225, 226, 233, 234, 242, 243, 261, 262, 269, 270, 278, 279, 297, 298, 305, 306, 314, 315, 333, 334, 341, 342, 350, 351, 369, 370, 371, 376, 377, 378, 379, 385, 386, 387, 406, 407, 408, 409, 410, 411, 412, 414, 415, 416, 420, 421, 422, 442, 443, 444, 445, 446, 447, 448, 450, 451, 452, 453, 454, 455, 456, 457, 458, 479, 480, 481, 482, 483, 487, 488, 489, 490, 491, 492, 493, 524, 525, 526, 527, 528:
					mask = 1;
				default: mask = 0;
			endcase
		end
		67: begin
			case(pos[9:0])
				51, 52, 53, 54, 55, 56, 57, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 155, 156, 157, 158, 166, 167, 168, 169, 170, 190, 191, 192, 204, 205, 206, 226, 227, 241, 242, 243, 261, 262, 263, 278, 279, 297, 298, 314, 315, 333, 334, 350, 351, 369, 370, 386, 387, 405, 406, 422, 423, 441, 442, 458, 459, 477, 478, 494, 495, 514, 515, 529, 530:
					mask = 1;
				default: mask = 0;
			endcase
		end
		68: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 206, 207, 225, 226, 242, 243, 261, 262, 278, 279, 297, 298, 314, 315, 333, 334, 350, 351, 369, 370, 371, 385, 386, 406, 407, 408, 420, 421, 422, 442, 443, 444, 445, 454, 455, 456, 457, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 554, 555, 556, 557, 558, 559, 560, 561:
					mask = 1;
				default: mask = 0;
			endcase
		end
		69: begin
			case(pos[9:0])
				117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 225, 226, 233, 234, 242, 243, 261, 262, 269, 270, 278, 279, 297, 298, 305, 306, 314, 315, 333, 334, 341, 342, 350, 351, 369, 370, 377, 378, 386, 387, 405, 406, 413, 414, 422, 423, 441, 442, 449, 450, 458, 459, 477, 478, 485, 486, 494, 495:
					mask = 1;
				default: mask = 0;
			endcase
		end
		70: begin
			case(pos[9:0])
				117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 225, 226, 234, 235, 261, 262, 270, 271, 297, 298, 306, 307, 333, 334, 342, 343, 369, 370, 378, 379, 405, 406, 414, 415, 441, 442, 450, 451, 477, 478, 486, 487:
					mask = 1;
				default: mask = 0;
			endcase
		end
		71: begin
			case(pos[9:0])
				51, 52, 53, 54, 55, 56, 57, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 155, 156, 157, 158, 166, 167, 168, 169, 170, 190, 191, 192, 204, 205, 206, 226, 227, 241, 242, 243, 261, 262, 263, 278, 279, 297, 298, 306, 307, 314, 315, 333, 334, 342, 343, 350, 351, 369, 370, 378, 379, 386, 387, 405, 406, 414, 415, 422, 423, 441, 442, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 477, 478, 486, 487, 488, 489, 490, 491, 492, 493, 494, 514, 515, 522, 523, 524, 525, 526, 527, 528, 529, 530:
					mask = 1;
				default: mask = 0;
			endcase
		end
		72: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 197, 198, 233, 234, 269, 270, 305, 306, 341, 342, 377, 378, 413, 414, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		73: begin
			case(pos[9:0])
				117, 118, 134, 135, 153, 154, 170, 171, 189, 190, 206, 207, 225, 226, 242, 243, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 369, 370, 386, 387, 405, 406, 422, 423, 441, 442, 458, 459, 477, 478, 494, 495:
					mask = 1;
				default: mask = 0;
			endcase
		end
		74: begin
			case(pos[9:0])
				117, 118, 133, 134, 153, 154, 170, 171, 189, 190, 206, 207, 225, 226, 242, 243, 261, 262, 278, 279, 297, 298, 314, 315, 333, 334, 349, 350, 351, 369, 370, 384, 385, 386, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492:
					mask = 1;
				default: mask = 0;
			endcase
		end
		75: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 198, 232, 233, 234, 235, 236, 267, 268, 269, 270, 271, 272, 273, 302, 303, 304, 307, 308, 309, 310, 336, 337, 338, 339, 345, 346, 347, 348, 371, 372, 373, 374, 382, 383, 384, 385, 406, 407, 408, 419, 420, 421, 422, 441, 442, 443, 457, 458, 459, 477, 478, 494, 495, 513, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		76: begin
			case(pos[9:0])
				117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 242, 243, 278, 279, 314, 315, 350, 351, 386, 387, 422, 423, 458, 459, 494, 495:
					mask = 1;
				default: mask = 0;
			endcase
		end
		77: begin
			case(pos[9:0])
				48, 49, 50, 51, 52, 53, 54, 55, 56, 57, 58, 59, 60, 61, 62, 63, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 191, 192, 193, 194, 195, 196, 230, 231, 232, 233, 234, 269, 270, 271, 272, 273, 307, 308, 309, 340, 341, 342, 343, 344, 372, 373, 374, 375, 376, 377, 405, 406, 407, 408, 409, 410, 441, 442, 443, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 560, 561, 562, 563, 564, 565, 566, 567:
					mask = 1;
				default: mask = 0;
			endcase
		end
		78: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 191, 192, 227, 228, 229, 230, 231, 265, 266, 267, 268, 269, 270, 304, 305, 306, 307, 308, 342, 343, 344, 345, 346, 347, 381, 382, 383, 384, 385, 420, 421, 422, 423, 441, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		79: begin
			case(pos[9:0])
				51, 52, 53, 54, 55, 56, 57, 58, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 154, 155, 156, 157, 158, 167, 168, 169, 170, 190, 191, 192, 205, 206, 207, 225, 226, 227, 241, 242, 243, 261, 262, 278, 279, 297, 298, 314, 315, 333, 334, 350, 351, 369, 370, 371, 385, 386, 387, 405, 406, 407, 420, 421, 422, 442, 443, 444, 445, 454, 455, 456, 457, 458, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 554, 555, 556, 557, 558, 559, 560, 561:
					mask = 1;
				default: mask = 0;
			endcase
		end
		80: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 199, 200, 225, 226, 235, 236, 261, 262, 271, 272, 297, 298, 307, 308, 333, 334, 343, 344, 369, 370, 371, 378, 379, 380, 406, 407, 408, 413, 414, 415, 442, 443, 444, 445, 446, 447, 448, 449, 450, 451, 479, 480, 481, 482, 483, 484, 485, 486, 516, 517, 518, 519, 520:
					mask = 1;
				default: mask = 0;
			endcase
		end
		81: begin
			case(pos[9:0])
				51, 52, 53, 54, 55, 56, 57, 58, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 154, 155, 156, 157, 158, 167, 168, 169, 170, 190, 191, 192, 205, 206, 207, 225, 226, 227, 241, 242, 243, 261, 262, 278, 279, 280, 281, 297, 298, 314, 315, 316, 317, 318, 319, 333, 334, 350, 351, 352, 353, 354, 355, 369, 370, 371, 385, 386, 387, 389, 390, 391, 392, 405, 406, 407, 420, 421, 422, 427, 428, 442, 443, 444, 445, 454, 455, 456, 457, 458, 463, 464, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 499, 500, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 535, 536, 554, 555, 556, 557, 558, 559, 560, 561, 570, 571, 572:
					mask = 1;
				default: mask = 0;
			endcase
		end
		82: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 99, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 189, 190, 197, 198, 225, 226, 233, 234, 261, 262, 269, 270, 297, 298, 305, 306, 307, 333, 334, 340, 341, 342, 343, 344, 369, 370, 371, 376, 377, 379, 380, 381, 382, 383, 406, 407, 408, 409, 410, 411, 412, 413, 416, 417, 418, 419, 420, 421, 422, 442, 443, 444, 445, 446, 447, 448, 454, 455, 456, 457, 458, 459, 480, 481, 482, 483, 493, 494, 495, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		83: begin
			case(pos[9:0])
				84, 85, 86, 87, 97, 98, 119, 120, 121, 122, 123, 124, 134, 154, 155, 156, 157, 158, 159, 160, 161, 170, 171, 190, 191, 195, 196, 197, 198, 206, 207, 225, 226, 227, 232, 233, 234, 242, 243, 261, 262, 269, 270, 278, 279, 297, 298, 305, 306, 307, 314, 315, 333, 334, 341, 342, 343, 350, 351, 369, 370, 378, 379, 380, 385, 386, 387, 405, 406, 414, 415, 416, 417, 421, 422, 441, 442, 451, 452, 453, 454, 455, 456, 457, 458, 478, 479, 487, 488, 489, 490, 491, 492, 493, 525, 526, 527, 528:
					mask = 1;
				default: mask = 0;
			endcase
		end
		84: begin
			case(pos[9:0])
				45, 46, 81, 82, 117, 118, 153, 154, 189, 190, 225, 226, 261, 262, 263, 264, 265, 266, 267, 268, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 297, 298, 299, 300, 301, 302, 303, 304, 305, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 369, 370, 405, 406, 441, 442, 477, 478, 513, 514, 549, 550:
					mask = 1;
				default: mask = 0;
			endcase
		end
		85: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 204, 205, 206, 241, 242, 243, 278, 279, 314, 315, 350, 351, 386, 387, 421, 422, 423, 456, 457, 458, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561, 562, 563:
					mask = 1;
				default: mask = 0;
			endcase
		end
		86: begin
			case(pos[9:0])
				45, 46, 47, 81, 82, 83, 84, 85, 86, 117, 118, 119, 120, 121, 122, 123, 124, 125, 156, 157, 158, 159, 160, 161, 162, 163, 164, 196, 197, 198, 199, 200, 201, 202, 203, 204, 235, 236, 237, 238, 239, 240, 241, 242, 243, 274, 275, 276, 277, 278, 279, 314, 315, 346, 347, 348, 349, 350, 351, 379, 380, 381, 382, 383, 384, 385, 386, 412, 413, 414, 415, 416, 417, 418, 419, 445, 446, 447, 448, 449, 450, 451, 452, 478, 479, 480, 481, 482, 483, 484, 485, 513, 514, 515, 516, 517, 518, 549, 550, 551:
					mask = 1;
				default: mask = 0;
			endcase
		end
		87: begin
			case(pos[9:0])
				81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 135, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 204, 205, 206, 207, 238, 239, 240, 241, 242, 243, 269, 270, 271, 272, 273, 274, 275, 276, 303, 304, 305, 339, 340, 341, 342, 343, 344, 345, 379, 380, 381, 382, 383, 384, 385, 418, 419, 420, 421, 422, 423, 457, 458, 459, 477, 478, 479, 480, 481, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 513, 514, 515, 516, 517, 518, 519, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531, 549, 550, 551, 552, 553, 554, 555, 556, 557, 558, 559, 560, 561:
					mask = 1;
				default: mask = 0;
			endcase
		end
		88: begin
			case(pos[9:0])
				27, 45, 62, 63, 81, 82, 96, 97, 98, 99, 117, 118, 119, 120, 131, 132, 133, 134, 135, 154, 155, 156, 157, 165, 166, 167, 168, 169, 191, 192, 193, 194, 195, 200, 201, 202, 203, 204, 228, 229, 230, 231, 232, 235, 236, 237, 238, 266, 267, 268, 269, 270, 271, 272, 273, 303, 304, 305, 306, 307, 338, 339, 340, 341, 342, 343, 344, 345, 373, 374, 375, 376, 378, 379, 380, 381, 382, 407, 408, 409, 410, 411, 416, 417, 418, 419, 420, 442, 443, 444, 445, 453, 454, 455, 456, 457, 477, 478, 479, 480, 491, 492, 493, 494, 495, 513, 514, 528, 529, 530, 531, 549, 566, 567:
					mask = 1;
				default: mask = 0;
			endcase
		end
		89: begin
			case(pos[9:0])
				9, 45, 46, 47, 81, 82, 83, 84, 118, 119, 120, 121, 122, 155, 156, 157, 158, 159, 160, 193, 194, 195, 196, 197, 231, 232, 233, 234, 235, 269, 270, 271, 272, 273, 274, 275, 276, 277, 278, 279, 306, 307, 308, 309, 310, 311, 312, 313, 314, 315, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 375, 376, 377, 378, 379, 409, 410, 411, 412, 413, 444, 445, 446, 447, 448, 478, 479, 480, 481, 482, 513, 514, 515, 516, 549, 550, 551:
					mask = 1;
				default: mask = 0;
			endcase
		end
		90: begin
			case(pos[9:0])
				81, 82, 98, 99, 117, 118, 133, 134, 135, 153, 154, 167, 168, 169, 170, 171, 189, 190, 201, 202, 203, 204, 205, 206, 207, 225, 226, 236, 237, 238, 239, 242, 243, 261, 262, 270, 271, 272, 273, 278, 279, 297, 298, 304, 305, 306, 307, 308, 314, 315, 333, 334, 339, 340, 341, 342, 350, 351, 369, 370, 373, 374, 375, 376, 386, 387, 405, 406, 407, 408, 409, 410, 411, 422, 423, 441, 442, 443, 444, 445, 458, 459, 477, 478, 479, 480, 494, 495, 513, 514, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		91: begin
			case(pos[9:0])
				151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 172, 173, 174, 175, 176, 177, 187, 188, 189, 190, 191, 192, 193, 194, 195, 196, 197, 198, 199, 200, 201, 202, 203, 204, 205, 206, 207, 208, 209, 210, 211, 212, 213, 223, 224, 225, 226, 227, 228, 229, 230, 231, 232, 233, 234, 235, 236, 237, 238, 239, 240, 241, 242, 243, 244, 245, 246, 247, 248, 249, 259, 260, 284, 285, 295, 296, 320, 321, 331, 332, 356, 357, 367, 368, 392, 393, 403, 404, 428, 429:
					mask = 1;
				default: mask = 0;
			endcase
		end
		92: begin
			case(pos[9:0])
				79, 115, 116, 117, 118, 151, 152, 153, 154, 155, 156, 190, 191, 192, 193, 194, 228, 229, 230, 231, 232, 233, 266, 267, 268, 269, 270, 271, 305, 306, 307, 308, 309, 310, 343, 344, 345, 346, 347, 348, 382, 383, 384, 385, 386, 420, 421, 422, 423, 424, 425, 458, 459, 460, 461, 462, 497, 498:
					mask = 1;
				default: mask = 0;
			endcase
		end
		93: begin
			case(pos[9:0])
				151, 152, 176, 177, 187, 188, 212, 213, 223, 224, 248, 249, 259, 260, 284, 285, 295, 296, 320, 321, 331, 332, 333, 334, 335, 336, 337, 338, 339, 340, 341, 342, 343, 344, 345, 346, 347, 348, 349, 350, 351, 352, 353, 354, 355, 356, 357, 367, 368, 369, 370, 371, 372, 373, 374, 375, 376, 377, 378, 379, 380, 381, 382, 383, 384, 385, 386, 387, 388, 389, 390, 391, 392, 393, 403, 404, 405, 406, 407, 408, 409, 410, 411, 412, 413, 414, 415, 416, 417, 418, 419, 420, 421, 422, 423, 424, 425, 426, 427, 428, 429:
					mask = 1;
				default: mask = 0;
			endcase
		end
		94: begin
			case(pos[9:0])
				124, 125, 158, 159, 160, 161, 193, 194, 195, 196, 197, 227, 228, 229, 230, 231, 261, 262, 263, 264, 297, 298, 333, 334, 335, 336, 370, 371, 372, 373, 408, 409, 410, 411, 445, 446, 447, 448, 449, 483, 484, 485, 520, 521:
					mask = 1;
				default: mask = 0;
			endcase
		end
		95: begin
			case(pos[9:0])
				32, 33, 68, 69, 104, 105, 140, 141, 176, 177, 212, 213, 248, 249, 284, 285, 320, 321, 356, 357, 392, 393, 428, 429, 464, 465, 500, 501, 536, 537, 572, 573:
					mask = 1;
				default: mask = 0;
			endcase
		end
		96: begin
			case(pos[9:0])
				151, 187, 188, 223, 224, 225, 259, 260, 261, 262, 296, 297, 298, 333, 334, 370:
					mask = 1;
				default: mask = 0;
			endcase
		end
		97: begin
			case(pos[9:0])
				94, 95, 96, 97, 122, 123, 128, 129, 130, 131, 132, 133, 134, 158, 159, 164, 165, 166, 167, 168, 169, 170, 171, 193, 194, 199, 200, 201, 205, 206, 207, 229, 230, 235, 236, 242, 243, 265, 266, 271, 272, 278, 279, 301, 302, 307, 308, 314, 315, 337, 338, 343, 344, 349, 350, 351, 373, 374, 379, 380, 385, 386, 409, 410, 411, 415, 416, 420, 421, 422, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 458, 459, 482, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 493, 494, 495, 520, 521, 522, 523, 524, 525, 526, 527, 528, 529, 530, 531:
					mask = 1;
				default: mask = 0;
			endcase
		end
		98: begin
			case(pos[9:0])
				79, 80, 81, 82, 83, 84, 85, 86, 87, 88, 89, 90, 91, 92, 93, 94, 95, 96, 97, 98, 115, 116, 117, 118, 119, 120, 121, 122, 123, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 134, 151, 152, 153, 154, 155, 156, 157, 158, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 171, 195, 196, 206, 207, 230, 231, 242, 243, 265, 266, 267, 278, 279, 301, 302, 314, 315, 337, 338, 350, 351, 373, 374, 385, 386, 387, 409, 410, 411, 412, 419, 420, 421, 422, 446, 447, 448, 449, 450, 451, 452, 453, 454, 455, 456, 457, 483, 484, 485, 486, 487, 488, 489, 490, 491, 492, 521, 522, 523, 524, 525, 526:
					mask = 1;
				default: mask = 0;
			endcase
		end
		99: begin
			case(pos[9:0])
				90, 91, 92, 93, 94, 95, 124, 125, 126, 127, 128, 129, 130, 131, 132, 133, 159, 160, 161, 162, 163, 164, 165, 166, 167, 168, 169, 170, 194, 195, 196, 197, 204, 205, 206, 229, 230, 231, 241, 242, 243, 265, 266, 278, 279, 301, 302, 314, 315, 337, 338, 350, 351, 373, 374, 386, 387, 409, 410, 422, 423, 446, 447, 457, 458:
					mask = 1;
				default: mask = 0;
			endcase
		end
		default: mask = 0;
	endcase
end

endmodule