`include "defines.v"

module rom(
	input wire[15:0] pc,
	output reg[15:0] ins_o
	);

	always @(*) begin
		//-*case*-/
		case (pc[15:0])
			16'h0000: ins_o = 16'b0110010000000000;    // MTSP R0
			16'h0001: ins_o = 16'b0000100000000000;    // NOP
			16'h0002: ins_o = 16'b0001000001000100;    // B START (START Addr=0x47)
			16'h0003: ins_o = 16'b0000100000000000;    // NOP
			16'h0004: ins_o = 16'b0000100000000000;    // NOP
			16'h0005: ins_o = 16'b0000100000000000;    // NOP
			16'h0006: ins_o = 16'b0000100000000000;    // NOP
			16'h0007: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0008: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0009: ins_o = 16'b0100111000010000;    // ADDIU R6 0x10
			16'h000a: ins_o = 16'b1101111000000000;    // SW R6 R0 0x00
			16'h000b: ins_o = 16'b1101111000100001;    // SW R6 R1 0x01
			16'h000c: ins_o = 16'b1101111001000010;    // SW R6 R2 0x02
			16'h000d: ins_o = 16'b1001000100000000;    // LW_SP R1 0x00
			16'h000e: ins_o = 16'b0110001100000001;    // ADDSP 0x01
			16'h000f: ins_o = 16'b0110100011111111;    // LI R0 0xFF
			16'h0010: ins_o = 16'b1110100100001100;    // AND R1 R0
			16'h0011: ins_o = 16'b1001001000000000;    // LW_SP R2 0x00
			16'h0012: ins_o = 16'b0110001100000001;    // ADDSP 0x01
			16'h0013: ins_o = 16'b0110001111111111;    // ADDSP 0xFF
			16'h0014: ins_o = 16'b1101001100000000;    // SW_SP R3 0x00
			16'h0015: ins_o = 16'b0110001111111111;    // ADDSP 0xFF
			16'h0016: ins_o = 16'b1101011100000000;    // SW_SP R7 0x00
			16'h0017: ins_o = 16'b0110101100001111;    // LI R3 0x0F
			16'h0018: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0019: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h001a: ins_o = 16'b0000100000000000;    // NOP
			16'h001b: ins_o = 16'b0001000010000001;    // B TESTW (TESTW Addr=0x9d)
			16'h001c: ins_o = 16'b0000100000000000;    // NOP
			16'h001d: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h001e: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h001f: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h0020: ins_o = 16'b0000100000000000;    // NOP
			16'h0021: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0022: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0023: ins_o = 16'b0000100000000000;    // NOP
			16'h0024: ins_o = 16'b0001000001111000;    // B TESTW (TESTW Addr=0x9d)
			16'h0025: ins_o = 16'b0000100000000000;    // NOP
			16'h0026: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0027: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0028: ins_o = 16'b1101111000100000;    // SW R6 R1 0x00
			16'h0029: ins_o = 16'b0000100000000000;    // NOP
			16'h002a: ins_o = 16'b0110101100001111;    // LI R3 0x0F
			16'h002b: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h002c: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h002d: ins_o = 16'b0000100000000000;    // NOP
			16'h002e: ins_o = 16'b0001000001101110;    // B TESTW (TESTW Addr=0x9d)
			16'h002f: ins_o = 16'b0000100000000000;    // NOP
			16'h0030: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0031: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0032: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h0033: ins_o = 16'b0000100000000000;    // NOP
			16'h0034: ins_o = 16'b0100001011000000;    // ADDIU3 R2 R6 0x00
			16'h0035: ins_o = 16'b1111001100000000;    // MFIH R3
			16'h0036: ins_o = 16'b0110100010000000;    // LI R0 0x80
			16'h0037: ins_o = 16'b0011000000000000;    // SLL R0 R0 0x0
			16'h0038: ins_o = 16'b1110101100001101;    // OR R3 R0
			16'h0039: ins_o = 16'b0110111110111111;    // LI R7 0xBF
			16'h003a: ins_o = 16'b0011011111100000;    // SLL R7 R7 0x00
			16'h003b: ins_o = 16'b0100111100010000;    // ADDIU R7 0x10
			16'h003c: ins_o = 16'b1001111100000000;    // LW R7 R0 0x00
			16'h003d: ins_o = 16'b1001111100100001;    // LW R7 R1 0x01
			16'h003e: ins_o = 16'b1001111101000010;    // LW R7 R2 0x02
			16'h003f: ins_o = 16'b1001011100000000;    // LW_SP R7 0x00
			16'h0040: ins_o = 16'b0110001100000001;    // ADDSP 0x01
			16'h0041: ins_o = 16'b0110001100000001;    // ADDSP 0x01
			16'h0042: ins_o = 16'b0000100000000000;    // NOP
			16'h0043: ins_o = 16'b1111001100000001;    // MTIH R3
			16'h0044: ins_o = 16'b1110111000000000;    // JR R6
			16'h0045: ins_o = 16'b1001001111111111;    // LW_SP R3 0xFF
			16'h0046: ins_o = 16'b0000100000000000;    // NOP
			16'h0047: ins_o = 16'b0110100000000111;    // LI R0 0x07
			16'h0048: ins_o = 16'b1111000000000001;    // MTIH R0
			16'h0049: ins_o = 16'b0110100010111111;    // LI R0 0xBF
			16'h004a: ins_o = 16'b0011000000000000;    // SLL R0 R0 0x00
			16'h004b: ins_o = 16'b0100100000010000;    // ADDIU R0 0x10
			16'h004c: ins_o = 16'b0110010000000000;    // MTSP R0
			16'h004d: ins_o = 16'b0000100000000000;    // NOP
			16'h004e: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h004f: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0050: ins_o = 16'b0100111000010000;    // ADDIU R6 0x10
			16'h0051: ins_o = 16'b0110100000000000;    // LI R0 0x00
			16'h0052: ins_o = 16'b1101111000000000;    // SW R6 R0 0x00
			16'h0053: ins_o = 16'b1101111000000001;    // SW R6 R0 0x01
			16'h0054: ins_o = 16'b1101111000000010;    // SW R6 R0 0x02
			16'h0055: ins_o = 16'b1101111000000011;    // SW R6 R0 0x03
			16'h0056: ins_o = 16'b1101111000000100;    // SW R6 R0 0x04
			16'h0057: ins_o = 16'b1101111000000101;    // SW R6 R0 0x05
			16'h0058: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0059: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h005a: ins_o = 16'b0000100000000000;    // NOP
			16'h005b: ins_o = 16'b0001000001000001;    // B TESTW (TESTW Addr=0x9d)
			16'h005c: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h005d: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h005e: ins_o = 16'b0110100001001111;    // LI R0 0x4F
			16'h005f: ins_o = 16'b1101111000000000;    // SW R6 R0 0x00
			16'h0060: ins_o = 16'b0000100000000000;    // NOP
			16'h0061: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0062: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0063: ins_o = 16'b0000100000000000;    // NOP
			16'h0064: ins_o = 16'b0001000000111000;    // B TESTW (TESTW Addr=0x9d)
			16'h0065: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0066: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0067: ins_o = 16'b0110100001001011;    // LI R0 0x4B
			16'h0068: ins_o = 16'b1101111000000000;    // SW R6 R0 0x00
			16'h0069: ins_o = 16'b0000100000000000;    // NOP
			16'h006a: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h006b: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h006c: ins_o = 16'b0000100000000000;    // NOP
			16'h006d: ins_o = 16'b0001000000101111;    // B TESTW (TESTW Addr=0x9d)
			16'h006e: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h006f: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0070: ins_o = 16'b0110100000001010;    // LI R0 0x0A
			16'h0071: ins_o = 16'b1101111000000000;    // SW R6 R0 0x00
			16'h0072: ins_o = 16'b0000100000000000;    // NOP
			16'h0073: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0074: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0075: ins_o = 16'b0000100000000000;    // NOP
			16'h0076: ins_o = 16'b0001000000100110;    // B TESTW (TESTW Addr=0x9d)
			16'h0077: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0078: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0079: ins_o = 16'b0110100000001101;    // LI R0 0x0D
			16'h007a: ins_o = 16'b1101111000000000;    // SW R6 R0 0x00
			16'h007b: ins_o = 16'b0000100000000000;    // NOP
			16'h007c: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h007d: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h007e: ins_o = 16'b0000100000000000;    // NOP
			16'h007f: ins_o = 16'b0001000000101000;    // B TESTR (TESTR Addr=0xa8)
			16'h0080: ins_o = 16'b0000100000000000;    // NOP
			16'h0081: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0082: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0083: ins_o = 16'b1001111000100000;    // LW R6 R1 0x00
			16'h0084: ins_o = 16'b0110111011111111;    // LI R6 0xff
			16'h0085: ins_o = 16'b1110100111001100;    // AND R1 R6
			16'h0086: ins_o = 16'b0000100000000000;    // NOP
			16'h0087: ins_o = 16'b0110100001010010;    // LI R0 0x52
			16'h0088: ins_o = 16'b1110100000101010;    // CMP R0 R1
			16'h0089: ins_o = 16'b0110000000110010;    // BTEQZ SHOWREGS (SHOWREGS Addr=0xbc)
			16'h008a: ins_o = 16'b0000100000000000;    // NOP
			16'h008b: ins_o = 16'b0110100001000100;    // LI R0 0x44
			16'h008c: ins_o = 16'b1110100000101010;    // CMP R0 R1
			16'h008d: ins_o = 16'b0110000001001101;    // BTEQZ SHOWMEM (SHOWMEM Addr=0xdb)
			16'h008e: ins_o = 16'b0000100000000000;    // NOP
			16'h008f: ins_o = 16'b0110100001000001;    // LI R0 0x41
			16'h0090: ins_o = 16'b1110100000101010;    // CMP R0 R1
			16'h0091: ins_o = 16'b0110000000100100;    // BTEQZ GOTOASM (GOTOASM Addr=0xb6)
			16'h0092: ins_o = 16'b0000100000000000;    // NOP
			16'h0093: ins_o = 16'b0110100001010101;    // LI R0 0x55
			16'h0094: ins_o = 16'b1110100000101010;    // CMP R0 R1
			16'h0095: ins_o = 16'b0110000000011101;    // BTEQZ GOTOUASM (GOTOUASM Addr=0xb3)
			16'h0096: ins_o = 16'b0000100000000000;    // NOP
			16'h0097: ins_o = 16'b0110100001000111;    // LI R0 0x47
			16'h0098: ins_o = 16'b1110100000101010;    // CMP R0 R1
			16'h0099: ins_o = 16'b0110000000011111;    // BTEQZ GOTOCOMPILE (GOTOCOMPILE Addr=0xb9)
			16'h009a: ins_o = 16'b0000100000000000;    // NOP
			16'h009b: ins_o = 16'b0001011111100000;    // B BEGIN (BEGIN Addr=0x7c)
			16'h009c: ins_o = 16'b0000100000000000;    // NOP
			16'h009d: ins_o = 16'b0000100000000000;    // NOP
			16'h009e: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h009f: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h00a0: ins_o = 16'b0100111000000001;    // ADDIU R6 0x01
			16'h00a1: ins_o = 16'b1001111000000000;    // LW R6 R0 0x00
			16'h00a2: ins_o = 16'b0110111000000001;    // LI R6 0x01
			16'h00a3: ins_o = 16'b1110100011001100;    // AND R0 R6
			16'h00a4: ins_o = 16'b0010000011111000;    // BEQZ R0 TESTW (TESTW Addr=0x9d)
			16'h00a5: ins_o = 16'b0000100000000000;    // NOP
			16'h00a6: ins_o = 16'b1110111100000000;    // JR R7
			16'h00a7: ins_o = 16'b0000100000000000;    // NOP
			16'h00a8: ins_o = 16'b0000100000000000;    // NOP
			16'h00a9: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h00aa: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h00ab: ins_o = 16'b0100111000000001;    // ADDIU R6 0x01
			16'h00ac: ins_o = 16'b1001111000000000;    // LW R6 R0 0x00
			16'h00ad: ins_o = 16'b0110111000000010;    // LI R6 0x02
			16'h00ae: ins_o = 16'b1110100011001100;    // AND R0 R6
			16'h00af: ins_o = 16'b0010000011111000;    // BEQZ R0 TESTR (TESTR Addr=0xa8)
			16'h00b0: ins_o = 16'b0000100000000000;    // NOP
			16'h00b1: ins_o = 16'b1110111100000000;    // JR R7
			16'h00b2: ins_o = 16'b0000100000000000;    // NOP
			16'h00b3: ins_o = 16'b0000100000000000;    // NOP
			16'h00b4: ins_o = 16'b0001000010101010;    // B UASM (UASM Addr=0x15f)
			16'h00b5: ins_o = 16'b0000100000000000;    // NOP
			16'h00b6: ins_o = 16'b0000100000000000;    // NOP
			16'h00b7: ins_o = 16'b0001000001101100;    // B ASM (ASM Addr=0x124)
			16'h00b8: ins_o = 16'b0000100000000000;    // NOP
			16'h00b9: ins_o = 16'b0000100000000000;    // NOP
			16'h00ba: ins_o = 16'b0001000011101101;    // B COMPILE (COMPILE Addr=0x1a8)
			16'h00bb: ins_o = 16'b0000100000000000;    // NOP
			16'h00bc: ins_o = 16'b0110100100000110;    // LI R1 0x06
			16'h00bd: ins_o = 16'b0110101000000110;    // LI R2 0x06
			16'h00be: ins_o = 16'b0110100010111111;    // LI R0  0xBF
			16'h00bf: ins_o = 16'b0011000000000000;    // SLL R0 R0 0x00
			16'h00c0: ins_o = 16'b0100100000010000;    // ADDIU R0 0x10
			16'h00c1: ins_o = 16'b1110001000101111;    // SUBU R2 R1 R3
			16'h00c2: ins_o = 16'b1110000001100001;    // ADDU R0 R3 R0
			16'h00c3: ins_o = 16'b1001100001100000;    // LW R0 R3 0x00
			16'h00c4: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h00c5: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h00c6: ins_o = 16'b0000100000000000;    // NOP
			16'h00c7: ins_o = 16'b0001011111010101;    // B TESTW (TESTW Addr=0x9d)
			16'h00c8: ins_o = 16'b0000100000000000;    // NOP
			16'h00c9: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h00ca: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h00cb: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h00cc: ins_o = 16'b0011001101100011;    // SRA R3 R3 0x00
			16'h00cd: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h00ce: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h00cf: ins_o = 16'b0000100000000000;    // NOP
			16'h00d0: ins_o = 16'b0001011111001100;    // B TESTW (TESTW Addr=0x9d)
			16'h00d1: ins_o = 16'b0000100000000000;    // NOP
			16'h00d2: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h00d3: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h00d4: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h00d5: ins_o = 16'b0100100111111111;    // ADDIU R1 0xFF
			16'h00d6: ins_o = 16'b0000100000000000;    // NOP
			16'h00d7: ins_o = 16'b0010100111100110;    // BNEZ R1 LOOP (LOOP Addr=0xbe)
			16'h00d8: ins_o = 16'b0000100000000000;    // NOP
			16'h00d9: ins_o = 16'b0001011110100010;    // B BEGIN (BEGIN Addr=0x7c)
			16'h00da: ins_o = 16'b0000100000000000;    // NOP
			16'h00db: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h00dc: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h00dd: ins_o = 16'b0000100000000000;    // NOP
			16'h00de: ins_o = 16'b0001011111001001;    // B TESTR (TESTR Addr=0xa8)
			16'h00df: ins_o = 16'b0000100000000000;    // NOP
			16'h00e0: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h00e1: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h00e2: ins_o = 16'b1001111010100000;    // LW R6 R5 0x00
			16'h00e3: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h00e4: ins_o = 16'b1110110111001100;    // AND R5 R6
			16'h00e5: ins_o = 16'b0000100000000000;    // NOP
			16'h00e6: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h00e7: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h00e8: ins_o = 16'b0000100000000000;    // NOP
			16'h00e9: ins_o = 16'b0001011110111110;    // B TESTR (TESTR Addr=0xa8)
			16'h00ea: ins_o = 16'b0000100000000000;    // NOP
			16'h00eb: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h00ec: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h00ed: ins_o = 16'b1001111000100000;    // LW R6 R1 0x00
			16'h00ee: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h00ef: ins_o = 16'b1110100111001100;    // AND R1 R6
			16'h00f0: ins_o = 16'b0000100000000000;    // NOP
			16'h00f1: ins_o = 16'b0011000100100000;    // SLL R1 R1 0x00
			16'h00f2: ins_o = 16'b1110100110101101;    // OR R1 R5
			16'h00f3: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h00f4: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h00f5: ins_o = 16'b0000100000000000;    // NOP
			16'h00f6: ins_o = 16'b0001011110110001;    // B TESTR (TESTR Addr=0xa8)
			16'h00f7: ins_o = 16'b0000100000000000;    // NOP
			16'h00f8: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h00f9: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h00fa: ins_o = 16'b1001111010100000;    // LW R6 R5 0x00
			16'h00fb: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h00fc: ins_o = 16'b1110110111001100;    // AND R5 R6
			16'h00fd: ins_o = 16'b0000100000000000;    // NOP
			16'h00fe: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h00ff: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0100: ins_o = 16'b0000100000000000;    // NOP
			16'h0101: ins_o = 16'b0001011110100110;    // B TESTR (TESTR Addr=0xa8)
			16'h0102: ins_o = 16'b0000100000000000;    // NOP
			16'h0103: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0104: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0105: ins_o = 16'b1001111001000000;    // LW R6 R2 0x00
			16'h0106: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h0107: ins_o = 16'b1110101011001100;    // AND R2 R6
			16'h0108: ins_o = 16'b0000100000000000;    // NOP
			16'h0109: ins_o = 16'b0011001001000000;    // SLL R2 R2 0x00
			16'h010a: ins_o = 16'b1110101010101101;    // OR R2 R5
			16'h010b: ins_o = 16'b1001100101100000;    // LW R1 R3 0x00
			16'h010c: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h010d: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h010e: ins_o = 16'b0000100000000000;    // NOP
			16'h010f: ins_o = 16'b0001011110001101;    // B TESTW (TESTW Addr=0x9d)
			16'h0110: ins_o = 16'b0000100000000000;    // NOP
			16'h0111: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0112: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0113: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h0114: ins_o = 16'b0011001101100011;    // SRA R3 R3 0x00
			16'h0115: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0116: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0117: ins_o = 16'b0000100000000000;    // NOP
			16'h0118: ins_o = 16'b0001011110000100;    // B TESTW (TESTW Addr=0x9d)
			16'h0119: ins_o = 16'b0000100000000000;    // NOP
			16'h011a: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h011b: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h011c: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h011d: ins_o = 16'b0100100100000001;    // ADDIU R1 0x01
			16'h011e: ins_o = 16'b0100101011111111;    // ADDIU R2 0xFF
			16'h011f: ins_o = 16'b0000100000000000;    // NOP
			16'h0120: ins_o = 16'b0010101011101010;    // BNEZ R2 MEMLOOP (MEMLOOP Addr=0x10b)
			16'h0121: ins_o = 16'b0000100000000000;    // NOP
			16'h0122: ins_o = 16'b0001011101011001;    // B BEGIN (BEGIN Addr=0x7c)
			16'h0123: ins_o = 16'b0000100000000000;    // NOP
			16'h0124: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0125: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0126: ins_o = 16'b0000100000000000;    // NOP
			16'h0127: ins_o = 16'b0001011110000000;    // B TESTR (TESTR Addr=0xa8)
			16'h0128: ins_o = 16'b0000100000000000;    // NOP
			16'h0129: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h012a: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h012b: ins_o = 16'b1001111010100000;    // LW R6 R5 0x00
			16'h012c: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h012d: ins_o = 16'b1110110111001100;    // AND R5 R6
			16'h012e: ins_o = 16'b0000100000000000;    // NOP
			16'h012f: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0130: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0131: ins_o = 16'b0000100000000000;    // NOP
			16'h0132: ins_o = 16'b0001011101110101;    // B TESTR (TESTR Addr=0xa8)
			16'h0133: ins_o = 16'b0000100000000000;    // NOP
			16'h0134: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0135: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0136: ins_o = 16'b1001111000100000;    // LW R6 R1 0x00
			16'h0137: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h0138: ins_o = 16'b1110100111001100;    // AND R1 R6
			16'h0139: ins_o = 16'b0000100000000000;    // NOP
			16'h013a: ins_o = 16'b0011000100100000;    // SLL R1 R1 0x00
			16'h013b: ins_o = 16'b1110100110101101;    // OR R1 R5
			16'h013c: ins_o = 16'b0110100000000000;    // LI R0 0x00
			16'h013d: ins_o = 16'b1110100000101010;    // CMP R0 R1
			16'h013e: ins_o = 16'b0110000000011101;    // BTEQZ GOTOBEGIN (GOTOBEGIN Addr=0x15c)
			16'h013f: ins_o = 16'b0000100000000000;    // NOP
			16'h0140: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0141: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0142: ins_o = 16'b0000100000000000;    // NOP
			16'h0143: ins_o = 16'b0001011101100100;    // B TESTR (TESTR Addr=0xa8)
			16'h0144: ins_o = 16'b0000100000000000;    // NOP
			16'h0145: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0146: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0147: ins_o = 16'b1001111010100000;    // LW R6 R5 0x00
			16'h0148: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h0149: ins_o = 16'b1110110111001100;    // AND R5 R6
			16'h014a: ins_o = 16'b0000100000000000;    // NOP
			16'h014b: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h014c: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h014d: ins_o = 16'b0000100000000000;    // NOP
			16'h014e: ins_o = 16'b0001011101011001;    // B TESTR (TESTR Addr=0xa8)
			16'h014f: ins_o = 16'b0000100000000000;    // NOP
			16'h0150: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0151: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0152: ins_o = 16'b1001111001000000;    // LW R6 R2 0x00
			16'h0153: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h0154: ins_o = 16'b1110101011001100;    // AND R2 R6
			16'h0155: ins_o = 16'b0000100000000000;    // NOP
			16'h0156: ins_o = 16'b0011001001000000;    // SLL R2 R2 0x00
			16'h0157: ins_o = 16'b1110101010101101;    // OR R2 R5
			16'h0158: ins_o = 16'b1101100101000000;    // SW R1 R2 0x00
			16'h0159: ins_o = 16'b0000100000000000;    // NOP
			16'h015a: ins_o = 16'b0001011111001001;    // B ASM (ASM Addr=0x124)
			16'h015b: ins_o = 16'b0000100000000000;    // NOP
			16'h015c: ins_o = 16'b0000100000000000;    // NOP
			16'h015d: ins_o = 16'b0001011100011110;    // B BEGIN (BEGIN Addr=0x7c)
			16'h015e: ins_o = 16'b0000100000000000;    // NOP
			16'h015f: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0160: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0161: ins_o = 16'b0000100000000000;    // NOP
			16'h0162: ins_o = 16'b0001011101000101;    // B TESTR (TESTR Addr=0xa8)
			16'h0163: ins_o = 16'b0000100000000000;    // NOP
			16'h0164: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0165: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0166: ins_o = 16'b1001111010100000;    // LW R6 R5 0x00
			16'h0167: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h0168: ins_o = 16'b1110110111001100;    // AND R5 R6
			16'h0169: ins_o = 16'b0000100000000000;    // NOP
			16'h016a: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h016b: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h016c: ins_o = 16'b0000100000000000;    // NOP
			16'h016d: ins_o = 16'b0001011100111010;    // B TESTR (TESTR Addr=0xa8)
			16'h016e: ins_o = 16'b0000100000000000;    // NOP
			16'h016f: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0170: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0171: ins_o = 16'b1001111000100000;    // LW R6 R1 0x00
			16'h0172: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h0173: ins_o = 16'b1110100111001100;    // AND R1 R6
			16'h0174: ins_o = 16'b0000100000000000;    // NOP
			16'h0175: ins_o = 16'b0011000100100000;    // SLL R1 R1 0x00
			16'h0176: ins_o = 16'b1110100110101101;    // OR R1 R5
			16'h0177: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0178: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0179: ins_o = 16'b0000100000000000;    // NOP
			16'h017a: ins_o = 16'b0001011100101101;    // B TESTR (TESTR Addr=0xa8)
			16'h017b: ins_o = 16'b0000100000000000;    // NOP
			16'h017c: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h017d: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h017e: ins_o = 16'b1001111010100000;    // LW R6 R5 0x00
			16'h017f: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h0180: ins_o = 16'b1110110111001100;    // AND R5 R6
			16'h0181: ins_o = 16'b0000100000000000;    // NOP
			16'h0182: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0183: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0184: ins_o = 16'b0000100000000000;    // NOP
			16'h0185: ins_o = 16'b0001011100100010;    // B TESTR (TESTR Addr=0xa8)
			16'h0186: ins_o = 16'b0000100000000000;    // NOP
			16'h0187: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0188: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0189: ins_o = 16'b1001111001000000;    // LW R6 R2 0x00
			16'h018a: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h018b: ins_o = 16'b1110101011001100;    // AND R2 R6
			16'h018c: ins_o = 16'b0000100000000000;    // NOP
			16'h018d: ins_o = 16'b0011001001000000;    // SLL R2 R2 0x00
			16'h018e: ins_o = 16'b1110101010101101;    // OR R2 R5
			16'h018f: ins_o = 16'b1001100101100000;    // LW R1 R3 0x00
			16'h0190: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h0191: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h0192: ins_o = 16'b0000100000000000;    // NOP
			16'h0193: ins_o = 16'b0001011100001001;    // B TESTW (TESTW Addr=0x9d)
			16'h0194: ins_o = 16'b0000100000000000;    // NOP
			16'h0195: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h0196: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h0197: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h0198: ins_o = 16'b0011001101100011;    // SRA R3 R3 0x00
			16'h0199: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h019a: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h019b: ins_o = 16'b0000100000000000;    // NOP
			16'h019c: ins_o = 16'b0001011100000000;    // B TESTW (TESTW Addr=0x9d)
			16'h019d: ins_o = 16'b0000100000000000;    // NOP
			16'h019e: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h019f: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h01a0: ins_o = 16'b1101111001100000;    // SW R6 R3 0x00
			16'h01a1: ins_o = 16'b0100100100000001;    // ADDIU R1 0x01
			16'h01a2: ins_o = 16'b0100101011111111;    // ADDIU R2 0xFF
			16'h01a3: ins_o = 16'b0000100000000000;    // NOP
			16'h01a4: ins_o = 16'b0010101011101010;    // BNEZ R2 UASMLOOP (UASMLOOP Addr=0x18f)
			16'h01a5: ins_o = 16'b0000100000000000;    // NOP
			16'h01a6: ins_o = 16'b0001011011010101;    // B BEGIN (BEGIN Addr=0x7c)
			16'h01a7: ins_o = 16'b0000100000000000;    // NOP
			16'h01a8: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h01a9: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h01aa: ins_o = 16'b0000100000000000;    // NOP
			16'h01ab: ins_o = 16'b0001011011111100;    // B TESTR (TESTR Addr=0xa8)
			16'h01ac: ins_o = 16'b0000100000000000;    // NOP
			16'h01ad: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h01ae: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h01af: ins_o = 16'b1001111010100000;    // LW R6 R5 0x00
			16'h01b0: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h01b1: ins_o = 16'b1110110111001100;    // AND R5 R6
			16'h01b2: ins_o = 16'b0000100000000000;    // NOP
			16'h01b3: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h01b4: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h01b5: ins_o = 16'b0000100000000000;    // NOP
			16'h01b6: ins_o = 16'b0001011011110001;    // B TESTR (TESTR Addr=0xa8)
			16'h01b7: ins_o = 16'b0000100000000000;    // NOP
			16'h01b8: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h01b9: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h01ba: ins_o = 16'b1001111001000000;    // LW R6 R2 0x00
			16'h01bb: ins_o = 16'b0110111011111111;    // LI R6 0xFF
			16'h01bc: ins_o = 16'b1110101011001100;    // AND R2 R6
			16'h01bd: ins_o = 16'b0000100000000000;    // NOP
			16'h01be: ins_o = 16'b0011001001000000;    // SLL R2 R2 0x00
			16'h01bf: ins_o = 16'b1110101010101101;    // OR R2 R5
			16'h01c0: ins_o = 16'b0100001011000000;    // ADDIU3 R2 R6 0x00
			16'h01c1: ins_o = 16'b0110111110111111;    // LI R7 0xBF
			16'h01c2: ins_o = 16'b0011011111100000;    // SLL R7 R7 0x00
			16'h01c3: ins_o = 16'b0100111100010000;    // ADDIU R7 0x10
			16'h01c4: ins_o = 16'b1001111110100101;    // LW R7 R5 0x05
			16'h01c5: ins_o = 16'b0110001111111111;    // ADDSP 0xFF
			16'h01c6: ins_o = 16'b1101010100000000;    // SW_SP R5 0x00
			16'h01c7: ins_o = 16'b1111010100000000;    // MFIH R5
			16'h01c8: ins_o = 16'b0110100110000000;    // LI R1 0x80
			16'h01c9: ins_o = 16'b0011000100100000;    // SLL R1 R1 0x0
			16'h01ca: ins_o = 16'b1110110100101101;    // OR R5 R1
			16'h01cb: ins_o = 16'b1001111100000000;    // LW R7 R0 0x00
			16'h01cc: ins_o = 16'b1001111100100001;    // LW R7 R1 0x01
			16'h01cd: ins_o = 16'b1001111101000010;    // LW R7 R2 0x02
			16'h01ce: ins_o = 16'b1001111101100011;    // LW R7 R3 0x03
			16'h01cf: ins_o = 16'b1001111110000100;    // LW R7 R4 0x04
			16'h01d0: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h01d1: ins_o = 16'b0100111100000100;    // ADDIU R7 0x04
			16'h01d2: ins_o = 16'b1111010100000001;    // MTIH R5
			16'h01d3: ins_o = 16'b1110111000000000;    // JR R6
			16'h01d4: ins_o = 16'b1001010100000000;    // LW_SP R5 0x00
			16'h01d5: ins_o = 16'b0000100000000000;    // NOP
			16'h01d6: ins_o = 16'b0000100000000000;    // NOP
			16'h01d7: ins_o = 16'b0110001100000001;    // ADDSP 0x01
			16'h01d8: ins_o = 16'b0110111110111111;    // LI R7 0xBF
			16'h01d9: ins_o = 16'b0011011111100000;    // SLL R7 R7 0x00
			16'h01da: ins_o = 16'b0100111100010000;    // ADDIU R7 0x10
			16'h01db: ins_o = 16'b1101111100000000;    // SW R7 R0 0x00
			16'h01dc: ins_o = 16'b1101111100100001;    // SW R7 R1 0x01
			16'h01dd: ins_o = 16'b1101111101000010;    // SW R7 R2 0x02
			16'h01de: ins_o = 16'b1101111101100011;    // SW R7 R3 0x03
			16'h01df: ins_o = 16'b1101111110000100;    // SW R7 R4 0x04
			16'h01e0: ins_o = 16'b1101111110100101;    // SW R7 R5 0x05
			16'h01e1: ins_o = 16'b1111000000000000;    // MFIH R0
			16'h01e2: ins_o = 16'b0110100101111111;    // LI R1 0x7F
			16'h01e3: ins_o = 16'b0011000100100000;    // SLL R1 R1 0x00
			16'h01e4: ins_o = 16'b0110101011111111;    // LI R2 0xFF
			16'h01e5: ins_o = 16'b1110100101001101;    // OR R1 R2
			16'h01e6: ins_o = 16'b1110100000101100;    // AND R0 R1
			16'h01e7: ins_o = 16'b1111000000000001;    // MTIH R0
			16'h01e8: ins_o = 16'b0110100100000111;    // LI R1 0x07
			16'h01e9: ins_o = 16'b1110111101000000;    // MFPC R7
			16'h01ea: ins_o = 16'b0100111100000011;    // ADDIU R7 0x03
			16'h01eb: ins_o = 16'b0000100000000000;    // NOP
			16'h01ec: ins_o = 16'b0001011010110000;    // B TESTW (TESTW Addr=0x9d)
			16'h01ed: ins_o = 16'b0000100000000000;    // NOP
			16'h01ee: ins_o = 16'b0110111010111111;    // LI R6 0xBF
			16'h01ef: ins_o = 16'b0011011011000000;    // SLL R6 R6 0x00
			16'h01f0: ins_o = 16'b1101111000100000;    // SW R6 R1 0x00
			16'h01f1: ins_o = 16'b0001011010001010;    // B BEGIN (BEGIN Addr=0x7c)
			16'h01f2: ins_o = 16'b0000100000000000;    // NOP
			default: ins_o = 16'h0800;
		endcase
		//-*case*-/
	end

endmodule